library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instr_mem is
    port(
        addr_instr : in std_logic_vector(31 downto 0);
        rd_instr : buffer std_logic_vector(31 downto 0)
    );
end instr_mem;

architecture rtl of instr_mem is

    type romtype is array (132 downto 0) of std_logic_vector(31 downto 0);
    signal mem : romtype;
     
begin
    
    -- mem(0) <= x"ff010113";
    -- mem(1) <= x"00812823";
    -- mem(2) <= x"01010413";
    -- mem(3) <= x"00400913";
    -- mem(4) <= x"ff242823";
    -- mem(5) <= x"00600913";
    -- mem(6) <= x"ff242a23";
    -- mem(7) <= x"00b00913";
    -- mem(8) <= x"ff242c23";
    -- mem(9) <= x"01100913";
    -- mem(10) <= x"ff242e23";
    -- mem(11) <= x"ffc42503";
    -- mem(12) <= x"ff842583";
    -- mem(13) <= x"ff840413";
    -- mem(14) <= x"00050463";
    -- mem(15) <= x"ff1ff0ef";
    -- mem(16) <= x"01010113";
    -- mem(17) <= x"00000013";
    -- mem(18) <= x"00000013";
    -- mem(19) <= x"00000013";
    -- mem(20) <= x"00000013";
    -- mem(21) <= x"00000013";
     mem(0)  <= x"ff010113";
     mem(1)  <= x"00812823";
     mem(2)  <= x"01010413";
     mem(3)  <= x"00400913";
     mem(4)  <=  x"ff242823";
     mem(5)  <= x"00600913";
     mem(6)  <= x"ff242a23";
     mem(7)  <=  x"00b00913";
     mem(8)  <= x"ff242c23";
     mem(9)  <= x"01100913";
     mem(10)  <= x"ff242e23";
     mem(11)  <= x"00000f13";
     mem(12)  <= x"ffc42503";
     mem(13)  <= x"ff842583";
     mem(14)  <= x"00000293";
     mem(15)  <= x"02300693";
     mem(16)  <= x"fff5c593";
     mem(17)  <= x"00b54533";
     mem(18)  <= x"00055e13";
     mem(19)  <= x"001e7393";
     mem(20)  <=  x"007282b3";
     mem(21)  <=  x"00155e13";
     mem(22)  <= x"001e7393";
     mem(23)  <= x"007282b3";
     mem(24)  <= x"00255e13";
     mem(25)  <= x"001e7393";
     mem(26)  <= x"007282b3";
     mem(27)  <= x"00355e13";
     mem(28)  <= x"001e7393";
     mem(29)  <= x"007282b3";
     mem(30)  <= x"00455e13";
     mem(31)  <= x"001e7393";
     mem(32)  <= x"007282b3";
     mem(33)  <=  x"00555e13";
     mem(34)  <= x"001e7393";
     mem(35)  <= x"007282b3";
     mem(36)  <= x"00655e13";
     mem(37)  <= x"001e7393";
     mem(38)  <= x"007282b3";
     mem(39)  <= x"00755e13";
     mem(40)  <= x"001e7393";
     mem(41)  <= x"007282b3";
     mem(42)  <= x"00855e13";
     mem(43)  <= x"001e7393";
     mem(44)  <= x"007282b3";
     mem(45)  <= x"00955e13";
     mem(46)  <= x"001e7393";
     mem(47)  <= x"007282b3";
     mem(48)  <= x"00a55e13";
     mem(49)  <= x"001e7393";
     mem(50)  <= x"007282b3";
     mem(51)  <= x"00b55e13";
     mem(52)  <= x"001e7393";
     mem(53)  <=  x"007282b3";
     mem(54)  <= x"00c55e13";
     mem(55)  <= x"001e7393";
     mem(56)  <= x"007282b3";
     mem(57)  <= x"00d55e13";
     mem(58)  <= x"001e7393";
     mem(59)  <=  x"007282b3";
     mem(60)  <= x"00e55e13";
     mem(61)  <= x"001e7393";
     mem(62)  <= x"007282b3";
     mem(63)  <= x"00f55e13";
     mem(64)  <=  x"001e7393";
     mem(65)  <= x"007282b3";
     mem(66)  <= x"01055e13";
     mem(67)  <= x"001e7393";
     mem(68)  <= x"007282b3";
     mem(69)  <= x"01155e13";
     mem(70)  <= x"001e7393";
     mem(71)  <= x"007282b3";
     mem(72)  <= x"01255e13";
     mem(73)  <= x"001e7393";
     mem(74)  <= x"007282b3";
     mem(75)  <= x"01355e13";
     mem(76)  <=  x"001e7393";
     mem(77)  <=  x"007282b3";
     mem(78)  <= x"01455e13";
     mem(79)  <=  x"001e7393";
     mem(80)  <= x"007282b3";
     mem(81)  <=  x"01555e13";
     mem(82)  <= x"001e7393";
     mem(83)  <=  x"007282b3";
     mem(84)  <=  x"01655e13";
     mem(85)  <=  x"001e7393";
     mem(86)  <= x"007282b3";
     mem(87)  <=  x"01755e13";
     mem(88)  <= x"001e7393";
     mem(89)  <=  x"007282b3";
     mem(90)  <=  x"01855e13";
     mem(91)  <=  x"001e7393";
     mem(92)  <=  x"007282b3";
     mem(93)  <=  x"01955e13";
     mem(94)  <= x"001e7393";
     mem(95)  <= x"007282b3";
     mem(96)  <= x"01a55e13";
     mem(97)  <=  x"001e7393";
     mem(98)  <= x"007282b3";
     mem(99)  <=  x"01b55e13";
     mem(100)  <= x"001e7393";
     mem(101)  <= x"007282b3";
     mem(102)  <= x"01c55e13";
     mem(103)  <= x"001e7393";
     mem(104)  <= x"007282b3";
     mem(105)  <= x"01d55e13";
     mem(106)  <= x"001e7393";
     mem(107)  <= x"007282b3";
     mem(108)  <= x"01e55e13";
     mem(109)  <= x"001e7393";
     mem(110)  <= x"007282b3";
     mem(111)  <= x"01f55e13";
     mem(112)  <= x"001e7393";
     mem(113)  <= x"007282b3";
     mem(114)  <= x"00500533";
     mem(115)  <= x"00151513";
     mem(116)  <= x"fe050293";
     mem(117)  <= x"005f0f33";
     mem(118)  <= x"00df4c63";
     mem(119)  <= x"00000013";
     mem(120)  <= x"00000013";
     mem(121)  <= x"00000013";
     mem(122)  <= x"00100e93";
     mem(123)  <= x"010000ef";
     mem(124)  <= x"00000e93";
     mem(125)  <= x"ff840413";
     mem(126)  <= x"e45ff0ef";
     mem(127)  <= x"01010113";
     mem(128)  <= x"00000013";
     mem(129)  <= x"00000013";
     mem(130)  <= x"00000013";
     mem(131)  <= x"00000013";
     mem(132)  <= x"00000013";

        process(addr_instr)begin
          rd_instr <= mem(to_integer(unsigned(addr_instr(31 downto 2))));
        end process;
    end rtl;
