library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity datapath is
    port(
        --inputs
        forward_ae      : in std_logic_vector(1 downto 0);
        forward_be      : in std_logic_vector(1 downto 0); 
        en_pc           : in std_logic;
        en_fd           : in std_logic;
        clr_fd          : in std_logic;
        clr_de          : in std_logic;
        clk             : in std_logic;
        reset           : in std_logic;
        pcsrc_e         : in std_logic;
        regwrite_d      : in std_logic;
        resultsrc_d     : in std_logic_vector(1 downto 0);
        memwrite_d      : in std_logic;
        jump_d          : in std_logic;
        branch_d        : in std_logic;
        alucontrol_d    : in std_logic_vector(2 downto 0);
        alusrc_d        : in std_logic;
        immsrc_d        : in std_logic_vector(1 downto 0);
        
        --outputs
        
        rd_e            : buffer std_logic_vector(4 downto 0);
        resultsrc_e     : buffer std_logic_vector(1 downto 0);
        regwrite_m      : buffer std_logic;
        rd_m            : buffer std_logic_vector(4 downto 0);
        rd_w            : buffer std_logic_vector(4 downto 0);
        instr_d         : buffer std_logic_vector(31 downto 0);
        zero_e          : out std_logic;
        jump_e          : out std_logic;
        branch_e        : out std_logic;
        rs1_e           : out std_logic_vector(4 downto 0);
        rs2_e           : out std_logic_vector(4 downto 0);
        regwrite_w      : buffer std_logic

    );
end datapath;

architecture rtl of datapath is

    --internal signals
    signal pcplus4_f        : std_logic_vector(31 downto 0);
    signal pcplus4_d        : std_logic_vector(31 downto 0);
    signal pctarget_e       : std_logic_vector(31 downto 0);
    signal pcf_in           : std_logic_vector(31 downto 0);
    signal pcf_buf          : std_logic_vector(31 downto 0);
    signal rd_instr         : std_logic_vector(31 downto 0);
    signal pc_d             : std_logic_vector(31 downto 0);
    signal rd_d             : std_logic_vector(4 downto 0);
    signal result_w         : std_logic_vector(31 downto 0);
    signal rd1              : std_logic_vector(31 downto 0);
    signal rd2              : std_logic_vector(31 downto 0);
    signal immext_d         : std_logic_vector(31 downto 0);
    signal regwrite_e       : std_logic;
    signal memwrite_e       : std_logic;
    signal alucontrol_e     : std_logic_vector(2 downto 0);
    signal alusrc_e         : std_logic;
    signal rd2_e            : std_logic_vector(31 downto 0);
    signal rd1_e            : std_logic_vector(31 downto 0);
    signal pc_e             : std_logic_vector(31 downto 0);
    signal immext_e         : std_logic_vector(31 downto 0);
    signal pcplus4_e        : std_logic_vector(31 downto 0);
    signal srcb_e           : std_logic_vector(31 downto 0);
    signal aluresult        : std_logic_vector(31 downto 0);
    signal writedata_e      : std_logic_vector(31 downto 0);      
    signal resultsrc_m      : std_logic_vector(1 downto 0);
    signal memwrite_m       : std_logic;
    signal aluresult_m      : std_logic_vector(31 downto 0);
    signal writedata_m      : std_logic_vector(31 downto 0);
    signal pcplus4_m        : std_logic_vector(31 downto 0);
    signal rd_memr          : std_logic_vector(31 downto 0);     
    signal resultsrc_w      : std_logic_vector(1 downto 0);
    signal aluresult_w      : std_logic_vector(31 downto 0);
    signal readdata_w       : std_logic_vector(31 downto 0);
    signal pcplus4_w        : std_logic_vector(31 downto 0);
    signal Src_AE           : std_logic_vector(31 downto 0);
    signal forward_be_mux_o : std_logic_vector(31 downto 0);
    
    
    begin
        --instantiation multiplexer 2 to 1
        inst_mux : entity work.mux_2(rtl)
            generic map(32)
            port map(
                port_in1    => pcplus4_f,
                port_in2    => pctarget_e,
                sel         => pcsrc_e,
                port_out    =>pcf_in
            );

        --instantiation program counter
        inst_pc : entity work.pc(rtl)
            port map(
                clk     => clk,
                reset   => reset,
                PCNext  => pcf_in,
                PC_cur  => pcf_buf,
                en      => en_pc 
            );

        --instantiation instruction memory
        inst_instr_mem : entity work.instr_mem(rtl)
            port map(
                addr_instr => pcf_buf,
                rd_instr => rd_instr
            );

        --instantiation adder +4
        inst_pcplus4 : entity work.PCPlus4(rtl)
            port map(
                a_in    => pcf_buf,
                b_in    => x"00000004",
                c_out   => pcplus4_f
            );

        --instantiation Register between fetch and decode
        inst_reg_fd : entity work.reg_fd(rtl)
            port map(
                clk         => clk,
                en          => en_fd,
                clr         => clr_fd,
                rd          => rd_instr,
                pc_f        => pcf_buf,
                pcplus4_f   => pcplus4_f,
                instr_d     => instr_d,
                pc_d        => pc_d,
                pcplus4_d   => pcplus4_d
            );

        --instantiation register file
        inst_reg_file : entity work.reg_file(rtl)
            port map(
                read_port_addr1     => instr_d(19 downto 15),
                read_port_addr2     => instr_d(24 downto 20),
                write_port_addr     => rd_w,
                write_data          => result_w,
                write_en            => regwrite_w,
                clk                 => clk,
                read_data1          => rd1,
                read_data2          => rd2
            );

        --instantiation extend
        inst_extend : entity work.extend(rtl)
            port map(
                ImmSrc => immsrc_d,
                instruction => instr_d(31 downto 7),
                ImmExt => immext_d
            );

        --instantiation Register between decode and execute
        inst_reg_de : entity work.reg_de(rtl)
            port map(
                clk             => clk,
                clr             => clr_de,
                regwrite_d      => regwrite_d,
                resultsrc_d     => resultsrc_d,
                memwrite_d      => memwrite_d,
                jump_d          => jump_d,
                branch_d        => branch_d,
                alucontrol_d    => alucontrol_d,
                alusrc_d        => alusrc_d,
                rd1             => rd1,
                rd2             => rd2,
                rs1_d           => instr_d(19 downto 15),
                rs2_d           => instr_d(24 downto 20),
                pc_d            => pc_d,
                rd_d            => rd_d,
                immext_d        => immext_d,
                pcplus4_d       => pcplus4_d,
                regwrite_e      => regwrite_e,
                resultsrc_e     => resultsrc_e,
                memwrite_e      => memwrite_e,
                jump_e          => jump_e,
                branch_e        => branch_e,
                alucontrol_e    => alucontrol_e,
                alusrc_e        => alusrc_e,
                rd1_e           => rd1_e,
                rd2_e           => rd2_e,
                rs1_e           => rs1_e,
                rs2_e           => rs2_e,
                pc_e            => pc_e,
                rd_e            => rd_e,
                immext_e        => immext_e,
                pcplus4_e       => pcplus4_e
            );

            
            --instantiation multiplexer 2 to 1
            inst_mux_2 : entity work.mux_2(rtl)
                generic map(32)
                port map(
                    port_in1    => forward_be_mux_o,
                    port_in2    => immext_e,
                    sel         => alusrc_e,
                    port_out    => srcb_e
                );
            
            --instantiation adder
            inst_adder : entity work.adder(rtl)
                port map(
                    a_in    => pc_e,
                    b_in    => immext_e,
                    c_out   => pctarget_e
                );
            
            --instantiation multiplexer for SrcAE
            inst_mux_3_src_ae : entity work.mux_3(rtl)
                generic map(32)
                port map(
                    port_in1    => rd1_e,
                    port_in2    => result_w,
                    port_in3    => aluresult_m,
                    sel         => forward_ae,
                    port_out    =>  Src_AE
                );
                
            --instantiation multiplexer for SrcBE
            inst_mux_3_src_be : entity work.mux_3(rtl)
                generic map(32)
                port map(
                    port_in1    => rd2_e,
                    port_in2    => result_w,
                    port_in3    => aluresult_m,
                    sel         => forward_be,
                    port_out    => forward_be_mux_o
                );
            --instantiation ALU
            inst_alu : entity work.ALU(rtl)
                port map(
                    SrcA            => Src_AE,
                    SrcB            => srcb_e,
                    ALUControl      => alucontrol_e,
                    Zero            => zero_e,
                    ALUResult       => aluresult
                );
            
            --instantiation Register between execute and memory
            writedata_e <= forward_be_mux_o;
            inst_reg_em : entity work.reg_em(rtl)
                port map(
                    clk             => clk,
                    regwrite_e      => regwrite_e,
                    resultsrc_e     => resultsrc_e,
                    memwrite_e      => memwrite_e,
                    aluresult       => aluresult,
                    writedata_e     => writedata_e,
                    rd_e            => rd_e,
                    pcplus4_e       => pcplus4_e,
                    regwrite_m      => regwrite_m,      
                    resultsrc_m     => resultsrc_m,
                    memwrite_m      => memwrite_m,
                    aluresult_m     => aluresult_m,
                    writedata_m     => writedata_m,
                    rd_m            => rd_m,
                    pcplus4_m       => pcplus4_m
                );

            --instantiation data memory
            inst_data_memr : entity work.data_memr(rtl)
                port map(
                    addr_port       => aluresult_m,
                    write_data      => writedata_m,
                    clk             => clk,
                    write_en        => memwrite_m,
                    read_data       => rd_memr
                );

            --instantiation Register between memory and writeback
            inst_reg_mw : entity work.reg_mw(rtl)
                port map(
                    clk             => clk,
                    regwrite_m      => regwrite_m,
                    resultsrc_m     => resultsrc_m,
                    aluresult_m     => aluresult_m,
                    rd              => rd_memr,
                    rd_m            => rd_m,
                    pcplus4_m       => pcplus4_m,
                    regwrite_w      => regwrite_w,    
                    resultsrc_w     => resultsrc_w,
                    aluresult_w     => aluresult_w,
                    readdata_w      => readdata_w,
                    rd_w            => rd_w,
                    pcplus4_w       => pcplus4_w
                );

            --instantiation multiplexer 3 to 1
            inst_mux_3 : entity work.mux_3(rtl)
                generic map(32)
                port map(
                    port_in1    => aluresult_w, 
                    port_in2    => readdata_w,
                    port_in3    => pcplus4_w,
                    sel         => resultsrc_w,
                    port_out    => result_w
                );
    end rtl;