library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instr_mem is
    port(
        addr_instr : in std_logic_vector(31 downto 0);
        rd_instr : buffer std_logic_vector(31 downto 0)
    );
end instr_mem;

architecture rtl of instr_mem is

    type romtype is array (135 downto 0) of std_logic_vector(31 downto 0);
    constant mem : romtype:=(
     x"ff010113",
     x"00812823",
     x"01010413",
     x"00400913",
     x"ff242823",
     x"00600913",
     x"ff242a23",
     x"00b00913",
     x"ff242c23",
     x"01100913",
     x"ff242e23",
     x"00000f13",
     x"ffc42503",
     x"ff842583",
     x"02000613",
     x"00000293",
     x"00000313",
     x"02300693",
     x"fff5c593",
     x"00b54533",
     x"00055e13",
     x"001e7393",
     x"007282b3",
     x"00155e13",
     x"001e7393",
     x"007282b3",
     x"00255e13",
     x"001e7393",
     x"007282b3",
     x"00355e13",
     x"001e7393",
     x"007282b3",
     x"00455e13",
     x"001e7393",
     x"007282b3",
     x"00555e13",
     x"001e7393",
     x"007282b3",
     x"00655e13",
     x"001e7393",
     x"007282b3",
     x"00755e13",
     x"001e7393",
     x"007282b3",
     x"00855e13",
     x"001e7393",
     x"007282b3",
     x"00955e13",
     x"001e7393",
     x"007282b3",
     x"00a55e13",
     x"001e7393",
     x"007282b3",
     x"00b55e13",
     x"001e7393",
     x"007282b3",
     x"00c55e13",
     x"001e7393",
     x"007282b3",
     x"00d55e13",
     x"001e7393",
     x"007282b3",
     x"00e55e13",
     x"001e7393",
     x"007282b3",
     x"00f55e13",
     x"001e7393",
     x"007282b3",
     x"01055e13",
     x"001e7393",
     x"007282b3",
     x"01155e13",
     x"001e7393",
     x"007282b3",
     x"01255e13",
     x"001e7393",
     x"007282b3",
     x"01355e13",
     x"001e7393",
     x"007282b3",
     x"01455e13",
     x"001e7393",
     x"007282b3",
     x"01555e13",
     x"001e7393",
     x"007282b3",
     x"01655e13",
     x"001e7393",
     x"007282b3",
     x"01755e13",
     x"001e7393",
     x"007282b3",
     x"01855e13",
     x"001e7393",
     x"007282b3",
     x"01955e13",
     x"001e7393",
     x"007282b3",
     x"01a55e13",
     x"001e7393",
     x"007282b3",
     x"01b55e13",
     x"001e7393",
     x"007282b3",
     x"01c55e13",
     x"001e7393",
     x"007282b3",
     x"01d55e13",
     x"001e7393",
     x"007282b3",
     x"01e55e13",
     x"001e7393",
     x"007282b3",
     x"01f55e13",
     x"001e7393",
     x"007282b3",
     x"00500533",
     x"00151513",
     x"fe050293",
     x"005f0f33",
     x"01e6d663",
     x"00300713",
     x"010000ef",
     x"00000e93",
     x"ff840413",
     x"e3dff0ef",
     x"01010113",
     x"00000013",
     x"00000013",
     x"00000013",
     x"00000013",
     x"00000013",
     x"00000013",
     x"00000013",
     x"00000013",
     x"00000013"
    );

    begin
    -- mem(136)    <= x"00000013";
    -- mem(137)    <= x"00000013";
    -- mem(138)    <= x"00000013";
    -- mem(139)    <= x"00000013";
    -- mem(140)    <= x"00000013";
        process(addr_instr)begin
          rd_instr <= mem(to_integer(unsigned(addr_instr(31 downto 0))));
        end process;
    end rtl;
